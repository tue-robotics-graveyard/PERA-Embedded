--------------------------------------------------------------------------------
-- Generated: 4-12-2014 15:06:40
--------------------------------------------------------------------------------
Library IEEE;
Use IEEE.Std_Logic_1164.all;
--------------------------------------------------------------------------------

--------------------------------------------------------------------------------
Entity Configurable_ADC_1 Is Port
--------------------------------------------------------------------------------
(
    DATA_I               : In   Std_Logic_Vector(15 DownTo 0);

    STB_I                : In   Std_Logic;
    CYC_I                : In   Std_Logic;
    ACK_O                : Out  Std_Logic;
    DAT_O                : Out  Std_Logic_Vector(15 DownTo 0);
    WE_I                 : In   Std_Logic;
    CLK_I                : In   Std_Logic;
    RST_I                : In   Std_Logic
);
--------------------------------------------------------------------------------
End Configurable_ADC_1;
--------------------------------------------------------------------------------

--------------------------------------------------------------------------------
Architecture Structure Of Configurable_ADC_1 Is
--------------------------------------------------------------------------------

    Signal IsReading                    : Std_Logic;
    Signal IsWriting                    : Std_Logic;
    Signal Acknowledge                  : Std_Logic;

    Signal ActiveAddress_DATA           : Std_Logic;

    Signal Read_DATA                    : Std_Logic;

--------------------------------------------------------------------------------
Begin
--------------------------------------------------------------------------------

    ----------------------------------------------------------------------------
    IsReading <= STB_I And CYC_I And Not WE_I;
    IsWriting <= STB_I And CYC_I And     WE_I;
    ----------------------------------------------------------------------------

    ----------------------------------------------------------------------------
    ACK_O <= Acknowledge;
    ----------------------------------------------------------------------------

    ----------------------------------------------------------------------------
    ActiveAddress_DATA <= '1';
    ----------------------------------------------------------------------------

    ----------------------------------------------------------------------------
    Process (IsReading, IsWriting, ActiveAddress_DATA)
    Begin
        Acknowledge      <= '0';
        Read_DATA        <= '0';

        If IsReading = '1' Then
            If ActiveAddress_DATA = '1'       Then Read_DATA <= '1';        Acknowledge  <= '1'; End If;
            If (ActiveAddress_DATA) = '0' Then Acknowledge <= '1'; End If;
        End If;
    End Process;
    ----------------------------------------------------------------------------

    ----------------------------------------------------------------------------
    Process (Read_DATA, DATA_I)
    Begin
        DAT_O <= (Others => '0');

        If Read_DATA = '1' Then
            DAT_O(15 DownTo 0) <= DATA_I;
        End If;
    End Process;
    ----------------------------------------------------------------------------

--------------------------------------------------------------------------------
End Structure;
--------------------------------------------------------------------------------
