library IEEE;
  use IEEE.std_logic_1164.all;
  use IEEE.numeric_std.all;

package adc_def is
  type adc_arr is array(0 to 7) of std_logic_vector(0 to 15);
end package adc_def;

