--------------------------------------------------------------------------------
-- Generated: 4-12-2014 15:06:40
--------------------------------------------------------------------------------
Library IEEE;
Use IEEE.Std_Logic_1164.all;
--------------------------------------------------------------------------------

--------------------------------------------------------------------------------
Entity Configurable_ENC_1 Is Port
--------------------------------------------------------------------------------
(
    C_I                  : In   Std_Logic_Vector(15 DownTo 0);

    STB_I                : In   Std_Logic;
    CYC_I                : In   Std_Logic;
    ACK_O                : Out  Std_Logic;
    DAT_O                : Out  Std_Logic_Vector(15 DownTo 0);
    WE_I                 : In   Std_Logic;
    CLK_I                : In   Std_Logic;
    RST_I                : In   Std_Logic
);
--------------------------------------------------------------------------------
End Configurable_ENC_1;
--------------------------------------------------------------------------------

--------------------------------------------------------------------------------
Architecture Structure Of Configurable_ENC_1 Is
--------------------------------------------------------------------------------

    Signal IsReading                    : Std_Logic;
    Signal IsWriting                    : Std_Logic;
    Signal Acknowledge                  : Std_Logic;

    Signal ActiveAddress_C              : Std_Logic;

    Signal Read_C                       : Std_Logic;

--------------------------------------------------------------------------------
Begin
--------------------------------------------------------------------------------

    ----------------------------------------------------------------------------
    IsReading <= STB_I And CYC_I And Not WE_I;
    IsWriting <= STB_I And CYC_I And     WE_I;
    ----------------------------------------------------------------------------

    ----------------------------------------------------------------------------
    ACK_O <= Acknowledge;
    ----------------------------------------------------------------------------

    ----------------------------------------------------------------------------
    ActiveAddress_C <= '1';
    ----------------------------------------------------------------------------

    ----------------------------------------------------------------------------
    Process (IsReading, IsWriting, ActiveAddress_C)
    Begin
        Acknowledge      <= '0';
        Read_C           <= '0';

        If IsReading = '1' Then
            If ActiveAddress_C = '1'          Then Read_C <= '1';           Acknowledge  <= '1'; End If;
            If (ActiveAddress_C) = '0' Then Acknowledge <= '1'; End If;
        End If;
    End Process;
    ----------------------------------------------------------------------------

    ----------------------------------------------------------------------------
    Process (Read_C, C_I)
    Begin
        DAT_O <= (Others => '0');

        If Read_C = '1' Then
            DAT_O(15 DownTo 0) <= C_I;
        End If;
    End Process;
    ----------------------------------------------------------------------------

--------------------------------------------------------------------------------
End Structure;
--------------------------------------------------------------------------------
